`define LOW       1'b0
`define HIGHT     1'b1

`define CMD_MODE  0
`define CMD_NOP   8
`define CMD_ANOP  24
`define CMD_ACTIV 3
`define CMD_WRITE 4
`define CMD_READ  5
`define CMD_PRECH 2

`define REG_MODE  12'h021

`define UNDEF32   32'bz
`define UNDEF16   16'bz